package pkg_msg;

parameter bit [7:0] POLY = 8'h9b;
parameter bit [7:0] BYTE_HEADER         = 8'h5a;
parameter bit [7:0] CMD_SINGLE_TRANS    = 8'hd1;

endpackage